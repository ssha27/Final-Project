module systolic_array(
    inp_west0,
    inp_west4,
    inp_west8,
    inp_west12,
    inp_north0,
    inp_north1,
    inp_north2,
    inp_north3,
    out00,
    out01,
    out02,
    out03,
    out04,
    out05,
    out06,
    out07,
    out08,
    out09,
    out10,
    out11,
    out12,
    out13,
    out14,
    out15,
	clk, 
    rst, 
    done);

// Your design is here




endmodule
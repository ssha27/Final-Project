

module PE(
    inp_north, 
    inp_west, 
    clk, 
    rst, 
    outp_south, 
    outp_east, 
    result);


// Your design is here

endmodule